package constants is
  constant DATA_WIDTH : natural := 32; -- bits
end package constants;