library IEEE;

use IEEE.std_logic_1164.all;
use WORK.tracker_constants.all;

entity i2c_tb is
end entity i2c_tb;

architecture behavioral of i2c_tb is

component i2c is
  generic (
    FREQUENCY : natural := 12_500_000 --10000
  );
  port (
    -- clocks
    clock_50 : in std_logic;
    reset : in std_logic;
    error : out std_logic;
    
    -- i2c communications
    sda : inout std_logic;
    scl : inout std_logic;
    data_clk : in std_logic;
    data_addr : in std_logic_vector(I2C_ADDR_WIDTH-1 downto 0);
    data_in : in std_logic_vector(I2C_DATA_WIDTH-1 downto 0);
    write_en, read_en : in std_logic; -- writing takes prescedence over reading
    available : out std_logic;
    
    -- fifo control
    write : in std_logic;
    odata : out std_logic_vector(7 downto 0);
    idata : in std_logic_vector(7 downto 0)
  );
end component i2c;

signal clock_50 : std_logic; --in
signal reset : std_logic; --in
signal error : std_logic; --out
signal sda : std_logic; --inout
signal scl : std_logic; --inout
signal data_clk : std_logic; --in
signal data_addr : std_logic_vector(I2C_ADDR_WIDTH-1 downto 0); --in
signal data_in : std_logic_vector(I2C_DATA_WIDTH-1 downto 0); --in
signal write_en : std_logic; --in
signal read_en : std_logic; --in
signal available : std_logic; --out
signal write : std_logic; --in
signal odata : std_logic_vector(7 downto 0); --out
signal idata : std_logic_vector(7 downto 0); --in
begin

test:i2c port map (clock_50, reset, error, sda, scl, data_clk, data_addr, data_in, write_en, read_en, available, write, odata, idata);

tester : process is
begin
	write_en <= '0';
	read_en <= '0';
	data_addr <= "1100011";
	data_in <= "11001100";
	
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	read_en <= '1';
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	read_en <= '0';
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	
	clock_50 <= '0';
	wait for 10 ns;
---------------------------------------------
	--sda <= '1';
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
--------------------------------------
	reset <= '1';
	write_en <= '1';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	reset <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;
	clock_50 <= '0';
	wait for 10 ns;
	clock_50 <= '1';
	wait for 10 ns;

wait;

end process tester;
end architecture behavioral;

